.title KiCad schematic
U1 Net-_R1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad2_ Net-_U1-Pad2_ Net-_C5-Pad2_ Net-_R1-Pad2_ Net-_R1-Pad2_ Net-_C4-Pad2_ Net-_R1-Pad2_ MAX256ASA
C4 Net-_C4-Pad1_ Net-_C4-Pad2_ C_Small
C5 Net-_C5-Pad1_ Net-_C5-Pad2_ C_Small
D3 Net-_C9-Pad2_ Net-_C4-Pad1_ Net-_C5-Pad1_ Net-_C9-Pad1_ D_Bridge_-AA+
D2 Net-_C4-Pad1_ Net-_C5-Pad1_ D_TVS
D1 Net-_C4-Pad2_ Net-_C5-Pad2_ D_TVS
C9 Net-_C9-Pad1_ Net-_C9-Pad2_ CP1
R1 Net-_R1-Pad1_ Net-_R1-Pad2_ R_Small
.end
